LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE work.components.all;

ENTITY InstructionMemory IS
    GENERIC(N : INTEGER := 32);
	PORT(
		Address				:IN STD_LOGIC_VECTOR ((N-1) DOWNTO 0);
		Instruction			:OUT STD_LOGIC_VECTOR ((N-1) DOWNTO 0)
		);
END InstructionMemory;

ARCHITECTURE Behavior OF InstructionMemory IS
BEGIN
 PROCESS(Address)
 BEGIN
    IF Address = "00000000000000000000000000000100" THEN
		Instruction <= "00001000000000010000000000000110"; -- addi R1,$ZERO,6 -> R1 <= 6
	ELSIF Address = "00000000000000000000000000001000" THEN
		Instruction <= "00001000000000100000000000001110"; -- addi R2,$ZERO,14 -> R2 <= 14
	ELSIF Address = "00000000000000000000000000001100" THEN
		Instruction <= "00001000000000110000000000001111"; -- addi R3,$ZERO,15 -> R3 <= 15
	ELSIF Address = "00000000000000000000000000010000" THEN
		Instruction <= "00001000000001000000000000011010"; -- addi R4,$ZERO,10 -> R4 <= 26
	ELSIF Address = "00000000000000000000000000010100" THEN
		Instruction <= "00001000000001010000000000001110"; -- addi R5,$ZERO,14 -> R5 <= 14
	ELSIF Address = "00000000000000000000000000011000" THEN
		Instruction <= "00001000000001100000000000100011"; -- addi R6,$ZERO,35 -> R6 <= 35
	ELSIF Address = "00000000000000000000000000011100" THEN
		Instruction <= "00001000000001110000000000010111"; -- addi R7,$ZERO,23 -> R7 <= 23
	ELSIF Address = "00000000000000000000000000100000" THEN
		Instruction <= "00001100010000100000000000000111"; -- subi R2,R2,7 => 14-7 = 7
	ELSIF Address = "00000000000000000000000000100100" THEN
		Instruction <= "00000000100001010010000000100010"; -- sub R4,R4,R5 => 26-14=12
	ELSIF Address = "00000000000000000000000000101000" THEN
		Instruction <= "00000000001001010001100000100000"; -- add R3,R1,R5 => 6+14=20
	ELSIF Address = "00000000000000000000000000101100" THEN
		Instruction <= "00000000110001010011000000100101"; -- or R6,R6,R5 => 35or14=47
	ELSIF Address = "00000000000000000000000000110000" THEN
		Instruction <= "00000000001000100000000000100100"; -- and R0,R1,R2 => 6and7=4
	ELSIF Address = "00000000000000000000000000110100" THEN
		Instruction <= "00001000101001010000000000000110"; -- addi R5,R5,6 -> R5 <= 6
	ELSIF Address = "00000000000000000000000000111000" THEN
		Instruction <= "00100100111000010000000000000011"; -- ori R1,R7,3 => 23or3=23
	ELSIF Address = "00000000000000000000000000111100" THEN
		Instruction <= "00011100011001100000000000000010"; -- andi R6,R3,2 => 20and2 = 2	
	ELSIF Address = "00000000000000000000000001000000" THEN
		Instruction <= "00010100010001000000000000000000"; -- sw R4,0(R2) => M7=12  
	ELSIF Address = "00000000000000000000000001000100" THEN
		Instruction <= "00110100000000000000000000000000"; -- NOP
	ELSIF Address = "00000000000000000000000001001000" THEN
		Instruction <= "00110100000000000000000000000000"; -- NOP
	ELSIF Address = "00000000000000000000000001001100" THEN
		Instruction <= "00101000101000110000000001000000"; -- beq R3,R5,BEQ(64)
	ELSIF Address = "00000000000000000000000001010000" THEN
		Instruction <= "00010000010000110000000000000000"; -- lw R3,0(R2)
	ELSIF Address = "00000000000000000000000001010100" THEN
		Instruction <= "00110100000000000000000000000000"; --NOP
	ELSE
		Instruction <= "00110100000000000000000000000000"; --NOP
  END IF;
 END PROCESS;
 
END Behavior;